library verilog;
use verilog.vl_types.all;
entity com_xnor_vlg_check_tst is
    port(
        ans_01          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end com_xnor_vlg_check_tst;
