library verilog;
use verilog.vl_types.all;
entity minu_time1_vlg_check_tst is
    port(
        CO_01           : in     vl_logic;
        Y_01            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end minu_time1_vlg_check_tst;
