library verilog;
use verilog.vl_types.all;
entity cnt12_vlg_vec_tst is
end cnt12_vlg_vec_tst;
