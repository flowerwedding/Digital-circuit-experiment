library verilog;
use verilog.vl_types.all;
entity Top_level_vlg_vec_tst is
end Top_level_vlg_vec_tst;
