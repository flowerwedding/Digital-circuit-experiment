library verilog;
use verilog.vl_types.all;
entity sys_choice_vlg_vec_tst is
end sys_choice_vlg_vec_tst;
