library verilog;
use verilog.vl_types.all;
entity bin_hour_vlg_vec_tst is
end bin_hour_vlg_vec_tst;
