library verilog;
use verilog.vl_types.all;
entity chron_vlg_vec_tst is
end chron_vlg_vec_tst;
