library verilog;
use verilog.vl_types.all;
entity minu_time1_vlg_vec_tst is
end minu_time1_vlg_vec_tst;
