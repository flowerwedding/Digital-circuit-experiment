library verilog;
use verilog.vl_types.all;
entity minu_time1_vlg_sample_tst is
    port(
        A0_01           : in     vl_logic;
        A1_01           : in     vl_logic;
        C1_01           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end minu_time1_vlg_sample_tst;
