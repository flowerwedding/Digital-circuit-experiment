library verilog;
use verilog.vl_types.all;
entity compare_vlg_check_tst is
    port(
        ans_01          : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end compare_vlg_check_tst;
