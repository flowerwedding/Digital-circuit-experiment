library verilog;
use verilog.vl_types.all;
entity m100 is
    port(
        pin_name2       : out    vl_logic;
        pin_name1       : in     vl_logic
    );
end m100;
