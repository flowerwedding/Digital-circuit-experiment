library verilog;
use verilog.vl_types.all;
entity minu_time1 is
    port(
        Y_01            : out    vl_logic;
        A0_01           : in     vl_logic;
        A1_01           : in     vl_logic;
        C1_01           : in     vl_logic;
        CO_01           : out    vl_logic
    );
end minu_time1;
