library verilog;
use verilog.vl_types.all;
entity bin_min_vlg_vec_tst is
end bin_min_vlg_vec_tst;
