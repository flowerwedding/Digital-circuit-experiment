library verilog;
use verilog.vl_types.all;
entity m100_vlg_check_tst is
    port(
        pin_name2       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end m100_vlg_check_tst;
