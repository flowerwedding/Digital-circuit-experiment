library verilog;
use verilog.vl_types.all;
entity minu60_vlg_vec_tst is
end minu60_vlg_vec_tst;
