library verilog;
use verilog.vl_types.all;
entity cnt100_vlg_vec_tst is
end cnt100_vlg_vec_tst;
