library verilog;
use verilog.vl_types.all;
entity seg_select_vlg_vec_tst is
end seg_select_vlg_vec_tst;
