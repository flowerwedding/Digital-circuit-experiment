library verilog;
use verilog.vl_types.all;
entity jicun_vlg_vec_tst is
end jicun_vlg_vec_tst;
