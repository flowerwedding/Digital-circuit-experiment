library verilog;
use verilog.vl_types.all;
entity bin_hour_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end bin_hour_vlg_sample_tst;
