library verilog;
use verilog.vl_types.all;
entity com_xnor_vlg_vec_tst is
end com_xnor_vlg_vec_tst;
