library verilog;
use verilog.vl_types.all;
entity chron_vlg_sample_tst is
    port(
        clk_01          : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end chron_vlg_sample_tst;
