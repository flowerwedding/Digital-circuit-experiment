library verilog;
use verilog.vl_types.all;
entity fre_div_vlg_vec_tst is
end fre_div_vlg_vec_tst;
