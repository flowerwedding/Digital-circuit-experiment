library verilog;
use verilog.vl_types.all;
entity minu60_vlg_sample_tst is
    port(
        clk_01          : in     vl_logic;
        CR_1            : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end minu60_vlg_sample_tst;
